interface dif;
	logic clk;
	logic rst_n;
	logic din;
	logic dout;
endinterface : dif